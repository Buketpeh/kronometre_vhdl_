library verilog;
use verilog.vl_types.all;
entity kronometreproje_vlg_vec_tst is
end kronometreproje_vlg_vec_tst;
